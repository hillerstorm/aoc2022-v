module days

fn test_day_eleven() {
	run_tests(day_eleven, [
		TestFixture{read_input(day: 11), '10605', '2713310158'},
	])
}
