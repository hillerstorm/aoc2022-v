module days

fn test_day_sixteen() {
	run_tests(day_sixteen, [
		TestFixture{read_input(day: 16), '1651', ''},
	])
}
