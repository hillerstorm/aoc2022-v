module days

fn test_day_thirteen() {
	run_tests(day_thirteen, [
		TestFixture{read_input(day: 13), '13', '140'},
	])
}
