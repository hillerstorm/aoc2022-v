module days

fn test_day_ten() {
	run_tests(day_ten, [
		TestFixture{read_input(day: 10), '13140', '
##..##..##..##..##..##..##..##..##..##..
###...###...###...###...###...###...###.
####....####....####....####....####....
#####.....#####.....#####.....#####.....
######......######......######......####
#######.......#######.......#######.....
'},
	])
}
