module days

fn test_day_seven() {
	run_tests(day_seven, [
		TestFixture{read_input(day: 7), '95437', '24933642'},
	])
}
