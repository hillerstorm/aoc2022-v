module days

fn test_day_fourteen() {
	run_tests(day_fourteen, [
		TestFixture{read_input(day: 14), '24', '93'},
	])
}
