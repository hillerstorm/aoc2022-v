module days

fn test_day_eight() {
	run_tests(day_eight, [
		TestFixture{read_input(day: 8), '21', '8'},
	])
}
